/* MODIFY. The cache controller. It is a state machine
that controls the behavior of the cache. */

module cache_control (
);

endmodule : cache_control
