module mp4();

endmodule : mp4
